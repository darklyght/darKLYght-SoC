module MMCMWrapper (
    output CLKFBOUT,
    output CLKFBOUTB,
    output CLKOUT0,
    output CLKOUT0B,
    output CLKOUT1,
    output CLKOUT1B,
    output CLKOUT2,
    output CLKOUT2B,
    output CLKOUT3,
    output CLKOUT3B,
    output CLKOUT4,
    output CLKOUT5,
    output CLKOUT6,
    input CLKFBIN,
    input CLKIN1,
    output LOCKED,
    input PWRDWN,
    input RST
);

    parameter BANDWIDTH = "OPTIMIZED",
              CLKOUT4_CASCADE = "FALSE",
              STARTUP_WAIT = "FALSE",
              CLKIN1_PERIOD = 0.000,
              DIVCLK_DIVIDE = 1,
              CLKFBOUT_MULT_F = 1.000,
              CLKFBOUT_PHASE = 0.000,
              CLKOUT0_DIVIDE_F = 1.000,
              CLKOUT0_PHASE = 0.000,
              CLKOUT0_DUTY_CYCLE = 0.500,
              CLKOUT1_DIVIDE = 1,
              CLKOUT1_PHASE = 0.000,
              CLKOUT1_DUTY_CYCLE = 0.500,
              CLKOUT2_DIVIDE = 1,
              CLKOUT2_PHASE = 0.000,
              CLKOUT2_DUTY_CYCLE = 0.500,
              CLKOUT3_DIVIDE = 1,
              CLKOUT3_PHASE = 0.000,
              CLKOUT3_DUTY_CYCLE = 0.500,
              CLKOUT4_DIVIDE = 1,
              CLKOUT4_PHASE = 0.000,
              CLKOUT4_DUTY_CYCLE = 0.500,
              CLKOUT5_DIVIDE = 1,
              CLKOUT5_PHASE = 0.000,
              CLKOUT5_DUTY_CYCLE = 0.500,
              CLKOUT6_DIVIDE = 1,
              CLKOUT6_PHASE = 0.000,
              CLKOUT6_DUTY_CYCLE = 0.500;

    MMCME2_BASE #(
        .BANDWIDTH(BANDWIDTH),
        .CLKOUT4_CASCADE(CLKOUT4_CASCADE),
        .STARTUP_WAIT(STARTUP_WAIT),
        .CLKIN1_PERIOD(CLKIN1_PERIOD),
        .DIVCLK_DIVIDE(DIVCLK_DIVIDE),
        .CLKFBOUT_MULT_F(CLKFBOUT_MULT_F),
        .CLKFBOUT_PHASE(CLKFBOUT_PHASE),
        .CLKOUT0_DIVIDE_F(CLKOUT0_DIVIDE_F),
        .CLKOUT0_PHASE(CLKOUT0_PHASE),
        .CLKOUT0_DUTY_CYCLE(CLKOUT0_DUTY_CYCLE),
        .CLKOUT1_DIVIDE(CLKOUT1_DIVIDE),
        .CLKOUT1_PHASE(CLKOUT1_PHASE),
        .CLKOUT1_DUTY_CYCLE(CLKOUT1_DUTY_CYCLE),
        .CLKOUT2_DIVIDE(CLKOUT2_DIVIDE),
        .CLKOUT2_PHASE(CLKOUT2_PHASE),
        .CLKOUT2_DUTY_CYCLE(CLKOUT2_DUTY_CYCLE),
        .CLKOUT3_DIVIDE(CLKOUT3_DIVIDE),
        .CLKOUT3_PHASE(CLKOUT3_PHASE),
        .CLKOUT3_DUTY_CYCLE(CLKOUT3_DUTY_CYCLE),
        .CLKOUT4_DIVIDE(CLKOUT4_DIVIDE),
        .CLKOUT4_PHASE(CLKOUT4_PHASE),
        .CLKOUT4_DUTY_CYCLE(CLKOUT4_DUTY_CYCLE),
        .CLKOUT5_DIVIDE(CLKOUT5_DIVIDE),
        .CLKOUT5_PHASE(CLKOUT5_PHASE),
        .CLKOUT5_DUTY_CYCLE(CLKOUT5_DUTY_CYCLE),
        .CLKOUT6_DIVIDE(CLKOUT6_DIVIDE),
        .CLKOUT6_PHASE(CLKOUT6_PHASE),
        .CLKOUT6_DUTY_CYCLE(CLKOUT6_DUTY_CYCLE)
    ) mmcm (
        .CLKFBOUT(CLKFBOUT),
        .CLKFBOUTB(CLKFBOUTB),
        .CLKOUT0(CLKOUT0),
        .CLKOUT0B(CLKOUT0B),
        .CLKOUT1(CLKOUT1),
        .CLKOUT1B(CLKOUT1B),
        .CLKOUT2(CLKOUT2),
        .CLKOUT2B(CLKOUT2B),
        .CLKOUT3(CLKOUT3),
        .CLKOUT3B(CLKOUT3B),
        .CLKOUT4(CLKOUT4),
        .CLKOUT5(CLKOUT5),
        .CLKOUT6(CLKOUT6),
        .CLKFBIN(CLKFBIN),
        .CLKIN1(CLKIN1),
        .LOCKED(LOCKED),
        .PWRDWN(PWRDWN),
        .RST(RST)
    );
    
endmodule
