 module OSERDESE2Wrapper #(
    parameter DATA_RATE_OQ = "DDR",
    parameter DATA_RATE_TQ = "DDR",
    parameter DATA_WIDTH = 1,
    parameter INIT_OQ = 1'b0,
    parameter INIT_TQ = 1'b0,
    parameter SERDES_MODE = "MASTER",
    parameter SRVAL_OQ = 1'b0,
    parameter SRVAL_TQ = 1'b0,
    parameter TBYTE_CTL = "FALSE",
    parameter TBYTE_SRC = "FALSE",
    parameter TRISTATE_WIDTH = 4
 ) (
    output OFB,
    output OQ,
    output SHIFTOUT1,
    output SHIFTOUT2,
    output TBYTEOUT,
    output TFB,
    output TQ,
    input CLK,
    input CLKDIV,
    input D1,
    input D2,
    input D3,
    input D4,
    input D5,
    input D6,
    input D7,
    input D8,
    input OCE,
    input RST,
    input SHIFTIN1,
    input SHIFTIN2,
    input T1,
    input T2,
    input T3,
    input T4,
    input TBYTEIN,
    input TCE
 );
    OSERDESE2 #(
        .DATA_RATE_OQ(DATA_RATE_OQ),
        .DATA_RATE_TQ(DATA_RATE_TQ),
        .DATA_WIDTH(DATA_WIDTH),
        .INIT_OQ(INIT_OQ),
        .INIT_TQ(INIT_TQ),
        .SERDES_MODE(SERDES_MODE),
        .SRVAL_OQ(SRVAL_OQ),
        .SRVAL_TQ(SRVAL_TQ),
        .TBYTE_CTL(TBYTE_CTL),
        .TBYTE_SRC(TBYTE_SRC),
        .TRISTATE_WIDTH(TRISTATE_WIDTH)
    ) oserdese2 (
        .OFB(OFB),
        .OQ(OQ),
        .SHIFTOUT1(SHIFTOUT1),
        .SHIFTOUT2(SHIFTOUT2),
        .TBYTEOUT(TBYTEOUT),
        .TFB(TFB),
        .TQ(TQ),
        .CLK(CLK),
        .CLKDIV(CLKDIV),
        .D1(D1),
        .D2(D2),
        .D3(D3),
        .D4(D4),
        .D5(D5),
        .D6(D6),
        .D7(D7),
        .D8(D8),
        .OCE(OCE),
        .RST(RST),
        .SHIFTIN1(SHIFTIN1),
        .SHIFTIN2(SHIFTIN2),
        .T1(T1),
        .T2(T2),
        .T3(T3),
        .T4(T4),
        .TBYTEIN(TBYTEIN),
        .TCE(TCE)
    );
    
endmodule
